���Uo� 3�3�?*N�fv�T���g�s�Q���Lno�R=FVu �Bq�եx�S���M����/f�NL�ܡ�Q�RO�=M.!)&}�y?�zŜx�R�xCS�"$0��̀�N�T��I���0���98�
^�䎐��!e)�9�����ӄla�q��I�q�ۺ!I	;�T�f�>�3��?d��z�O8y�̙�z
y�sAn�� �����d�������	0	�����k��Q�q�c�}}i�<�Pc���}� �z�2�\n#�x��܆3��h/�,D���ju��Eo�1�Kc�Ӝ�R-̌�f����
��Ph�Wrt�؟A�ә�}�?��t����]
X�w4�˳nd����~NV�Mn��Ȁό.6Ԓs��W�`82��r0~�.�E��<n�prG�5��`x�O���{����%�e�m�s��z���7����?1�� ������R���ĭ��e�f��8V��W�c��]}�O ��Uɵ��'��K� �4�!�a�qI� ��K��M�� ���� /��Rv�k�ɻb6c��?Z���~g�3�?:r��`����Ǳ.�$W��.����~��� �U��.3�O�s�����~i� ���S[�,>S�4}U�1�s1��dr6��W[�Dl��={{u�8*� 3���Q�:{�K�A�YQ�s+|��w���q���������ߊwq�:P��^�cg�c�<�V|