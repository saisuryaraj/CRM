M��Dr$���+ڼ5�x~M
�-݈�#$�_��~Q&��y�Ǭݿ#�N:zu�G���Z���ܲ��rߦ8���3�2��?J�`���I�X����lv�x��+�;���Kq-ǔ�1��?����F�>+��o�ۗ�8i?�?*٨�r=�D{6��Y�~
�!���閖[9m(s'n��yg�,M}Roc��1 �s�c��WEk���<�<�� �NI � �	�%��;����|ZCL`�c���rz�;֗ssIu �$t����>�����q�X]�2���9V$o�,�����PVI�Ѥћ��[ɥ��G3[H �����w��x�T���1}��Y0:s��1�����mJ��۝��T.[?�?�xַ�������r��d*	�돥\d>�U��\j,�N���Î3��=?
ߍn���E��إ�I��O#��� >6���$����Ʌ &��c��x=*�~
���q�R��ϧ^�ޕw3���\]����HZE� J�L0<��sW�.<Oi�i�isKÜ��	��ާ�>�7���?��I`rL��F<0�oa���^�yeb��Yۜi�Q�w{b���yg���;��2��y���GZ�״����#^�go�RxB!k��/�̜���:Wg�J��d�n�����q@��<�R���w��F�׍ǁ��ry�bi�Uŭ��8����������O���)#1a��d���k�Z��l��4�������XynpzⰯ�Z�hd��B6�$1�� �w�$�/.b2.Yʅl 9�W6�Z�S2䱌�FH������^ǔXM��>�WN��1���s�����z������$�T)۸8���k�ѓD��4H�"�HQ^1���OL��^��0�3��&L@q!A��T�a�8i�<��Q�L�ePU�9�Nk�{Yt�.��R�gհ2MqVs�C�^S4p���ҽ^��;��F4p�-�_����>��z�j~�V����~/�+]���>Qq� �oJ�&u��v�.�vc{�<��O�y�W��xZ���Ry4�)�]�y�qǾk��τ�,�"ڈ��J]nO��8�=�U▅YX�K�Q�2ݴἸ�6��װ��]�iر<���B�|�c��Y�-���.�~���0G�����_S�Ɨ�5�Pj.6��� �Ϛ��	�s������#�Xٷ�	���x%���$�l�k�JǑ�z���W�x���u8�,���LWB��X�sӡ=k˴=6�<m$v��(�3��V�D$���/��m�)�2jЫ-�$��I�;��#��L��K��׮q���u���������-���dd���b_x��S��^�3���ظ^rSY$��}L9�Akm�9}r��hN׍N�ݻg�i�4�k�/���*䜱'��Qkj�櫧�dG�|�!��8��g޵ZOi�?u��FS4*��NI�Zv@���v�>��X� ���.V @ �>���S���V7	>��;9��Y����0#�,�lr2N9��&��aY.�`W�"�V04�S\���4ԧ*˂�1 ���#����qf�\c���R՟Nf�B�=?�Yܫ�}���q��zT� �W8{�����ɿ� �:��ҦՄ��kw��qć�Zך��