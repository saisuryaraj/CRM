dZ��V����
��6}9��[/�t�(�x�=��W"�l��d�c��g�� �|Yk�
E*�'Ps�����b_j���2�nQ���	�ų��aI���$*��v�'���C� ��^�?Ӥ=�<�n�x�SH�s���� �Zd�3�ɵKmʿ'Ld�4K�em@M|�a��t̸m�7
��Jf�� B5JWbq�=�M���B���v>��N?��1�����Hs�+�(�l�|�'ߊ� l��Zq�3����H�3q�y� �V�̠�|��֫�`��>B7�ʹ�L��xnK-"# �;�j�iFҡ���ޛ:���y�I#��<f�|In������� �.f�$W��fO0�^O��Zv+�&�ݷ9#=�el���RQg��
�n��,x^{���v9lX�~�v:zU�J�G�隯6�����V�J<����V��j�z������)�s�g� �I���9=8�,09=x�cC@�8�NO��H��0S�N��~v�����6cvT|ǥFG�v5����C���@ɔ(���r;Tl�61���y�ߍB'����8w���g�֣����S�������\�1�T*A*rzԫ�~f�	0?N�*ݷ�cP��� ��S��(�:�I��%v/N�3N��{�F3'��?+���R�c<v�``���Ҥ�<��/ˎ߈�����w)S��^ߍ?��`�4�S�����"E8�i~� a�}�n�H?0� >�1r <�I&>���T�;~�S�����hD����B ���zՐ͐8�ґ���1�Vއ�4����1�>�Q��	?68�I�#s��U%a�I�Ǘ�5i�'��T&#ʘ��i�|�A6d�p��̜l��9�y�+����ӧoz�5'?j�Ỏ?
@q��Zy>��� j���>f8�Z�x@y�n�=���o�H���G��,�
Ǌ�|���ua�e���^q�p~�o���J�'��m�Խ��Ǩ� ��z�`��v���j�v/�L��Q2� ����ַ�� ��_�+
<y��[��d��ҹ�n�m_?�����E|�㹁�QU�����^u�%��f��'���_�)� X~��皠�ؔ{�iZ��Q�gNǀj�x�r3W�������;-?>m��+�t��L
Kt�t�>��{V/A��Oʻ�6�l�~z���GQ�8O���a�˭h�ؕ9^������
I��|9ll�l��(�$m��V�W�k63��c��*��ÓT�.�e�#�� �V#c��֩.B� ���H~O��S}s�ӗ93u5l0����e6�v�	�,p:ӕ�' ����h c��1x�=H���j�ױ�&2x;P&X��JU�y��h�:�R�BW��q$J'�c'�J���T��ǃ��2�-�qHe�~Sӯz� ��1�Ԝ���A���h&x�)	�������:Sn�8��4�=s׽
~q��QH��3`E�*z��2`W'�N�hS��T���� ;��c���N@2� �۵JTn&�0i��� o�(�( y�*�%!��O'��39#�8�1��}�
�l�8���J�D#��_�~��i�>\q�T�x�>�+s��u�i���4�>n�����6x�����*��PH8jLh�b|�庚�\���i
�x?z��8l`T�X�>�T��<�+T� �G���L��P���N��x<�J���X�囯�IC��z���t=;T�`�^i��'ʡ���\�G=�0�1�D$ �0���!;׭C�p[�X��� j�iSx��:H���o�J�&Y\�^��Fx��D�#�5f2w��1�W<�J�P�w=�z�' o���Sb����?z�O���t����3}�ɕ�$d�R�K��-�k<��ס��8�[��TX���қ7'ʓ��;�)'�u�bs���9�B��q��s�h��c����k9+3zN���1�0|a��d(��T}A5�60y��98��^��^�!�ѭH�5��(���s^G*1G
8kX�V'�*����~���pNޤ(�