�l`{��y�#��7þ#��[����H8�u�ς�+k�6}0mU��}3�Ƶ��a̡��z]���񉴬�A�%�������/P1]Wbd�:c����Ƒ����6x^�m|9l�d����c�j�TÞ�v���nˣ�J��� �ҵ������B/���ٓ�s_X���7���m� g��g���m������*���>#��]�g?غ���C�������j����ԉ�1�dҿA'�f����m����.����f�Н�N�I�j��畍������5Dh�#=x'���}E�_:��A��>~����^�k�+��ߞk:/\D\G-��}r,�~�,�(x���?��[$����9�Ex%���g�#��ۼ}���Lq�8���M��W�Ksd� y�??��w_������������48NV>f�5Sif�3�'�>��r?�I!��K~�p?¾��𞔥G�&���D:U��=�� �5���STE� |��⹕cm2��K�~Q����5�W�� �G���k쨼3������� @��8=�hg?�,�|��y�������O֞ �A��� ���*�[��˧jck��C�ȁ_j� �?��`t�b3�?�R�Ь�D�h�{ Dgc���h�?}�(�8��>ai���8�;W�?�X��8�,ă��?Z�?��3i���aܥ�E`:v {����+���ggwɐ�H�W#vf�Χ�����-�RrOr}}�^���~֤q¾GҼC���Y$22UP�p�J�}�K�H�il'	�W����i�L繢�3i2���-��Es:����2)0�һ&���}ҟ�������F�Mr��Axa����`�c�4�8��<^]����֓����Wf��c��� 'j�z������M/n���s�>��;���qF7��u�O�\1��Q�W֟�=OZ1}:S�N���Fr)�u�h���iy�Ґ���;R��@�^���zA�OJ^7u4 ��Q����:u�u�җ��@�ۥ ��;��h;��O�?x�� �����i ��OΎǯZ_^E�ҕ�`�G�)pq׵4�'���`����0��?.7zR���i��2}i�F����9ǽE�erǿ~��iTzJ���e��Q�í ͙��vS$A���a�_�������^� �s��I%��쇑���BI�/�&	��$Ӓ�������;�a����=�����C��<g�z�϶.ܑ�@�a�n��è�rG��*2Ҏ�N� $������@D���nǷ>�;�N���s�{gڠc�-�%�9n����Tʤ���#5eW��x�#`4X\�C���#� �I�����6�$c���P!/�N��껲���#������f?^�ӎ��Xc�ز����#�� �PH���U���L�3ݺ��T�H�A��@K���A������c==G�W�.m�\c�+7;�PI��z㿵4��Y��?pw��V��y�Q1��X�����'��������Z��"��f�F����Mzlg�ɼ���q_\h�Ů�l�d،p�� Z���;K	iʶ�Z���	@� u�����S�6�9�-���UҴ������į�zMލ�\[�vv��D��