�Xw8xt����G=GlՔ�6����PG<?*�J��qC�&��c;�.FW;N:��N䘑X"��c�+Eb�܎���U�X����<�g͸����� �ZN�Ҟq��zO_��Bhi�w���ގ�i�C��L�/��c��t�aӃ�֐���J1�޴�1ӵ(ϥ��1�=������!�7j��?4���z�J\�9��>��!�9�Vt���~�À1��U�K.ӵt�E���[�h���������O	 ��1%��@��a]���j�z|��^?1�ָ=&'�MM�6��>P��O��H���BO� ������z����-�9�����*kӂH��^���\�$cV�-��� �u7��-�,��`�>�Q�\\�}�j�;ˍ��v� ?J��߈"ٛ�)��py�=��Y�߇v�q'C��]���6q�O��z
���<����r>\�������m-��͟���^}ogp��|��2�9?��W�k�z" �$�#=��AӚk�w{C��X珥�S�:/@V�" ~cR�5)�;��w�O5�Z[���I�����+��l�R �?9�c�_)�w0���B{��������7*`�>�A�d��2�p0k1o'���	���Jm	�};ọ:;!�y_���[��E�G�c��|��k�F�7�b{���ؚ�;V���b� .�p=?�j!&��n�c���|�� %^3�������F����s���������t`?���Z�ս�Ω�|»��|�-A�Q�!����8��v� *��LwX��˂;k�i�A#/�b�޷t�Ke�"=�&��=MK�&���.�s�2C�c�� J���*K{�]�2��z��S��r�Z?ƼGŶ�4�q�,�`z�?��qL�2����t7�.��m#�#�zU��maW�$W�� *�|5mq&�jM�W�x�^�>��M��0<���?�e*Z�9�����Q�:�k6H]B�}�݉�|̼�[���P�� ���Cu!�����Y�w��Q��b4�H��������i�1lc��?�u6�7+��ܑ�z��_G�2�(A����ǰ{Yc���Ƥ���l��T㽃�����D�~��|D��m7�ϝ�XW�>+��v�f,=�F'Tj;z\~����|p}����җ���B��}��t� 0�!%�9�3��5*�>W��£�.��Fo�2\͸�d2g ������9���Y�tOg�?�*_� #3|:^�;5#�aɐ��Ҕ�f�ڧ�EV�BƳ~�	��� �����ޞ�H[�X�#`d�;u��!��+5���� hK��ha��i$�zO�'����0'Ձ��1�}jQ4%]�yX'<�ڡ��b�fk4��!��S�g.z�^3�)������\���z�� �V�-���?Ձ���΄ts�q�Q�e�~ݚFF)�qʢ�O9��8\^"��<��O�f��oC��9�?̈$K����K��?�2��Nc)�p�c�E��!��6XAǥSA���1��� �z�|!s�do?\R��{�e�#3�N������S��\X����A�̿�`��R����G0��#����.�*���t�I�����O� �1��8ϯ|V+c#3�y�
����cn~`ϯ�f�Qn����Ȫ�ۈ�z~��.E;y��X�y��r����z�g?6\��1O�q�/n�tĺmjO��69����*7sT@>c}���H�$���Z_R]���o��62��I*yoaY�N˨����ߝU�~_M��TNْ>8�j��!�`֚�h��9��� ֨b�,�N6	�`o������ `������(=�zY�:r=�Ҷb�b@{n{o��a�
2�1�K�N�,nG��pD� ��D�e*��2�rg,>ҿ�ӟ�]	�AR�H���9� 
�C�F� Y̹�?���