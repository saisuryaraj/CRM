y=9�/c��)��s~=s�LL�E��eOL�U#m'�N�s�*�<7#�0� �?1�rGY��`��� _T�8���â�i�~A��ׯZ�aFUpː8�v���c-��:�9`L�� �"̪ŵ��ܺo�����=p�<F��b�4h��Xi�Ir�y���x��|m.�6j�l|���q��j�x��-!-=�>x��P � �U_��F]ϫb�I6�d�r�r '׏�W�z_��f����_*��<\"R5{�å9�Q�a��ڎ��2W��|���>�J��ش�pR	�;��^�<���u�q����I�o��n����J�� 	G�Xs��_�o��M? �����k`�l,:s�rER�Z��V;,��qbz��m߉|Z�E[T��A'� �+:�]��m�=N��C��׏���3�%M5��w	�LU;�m���h,@c�������Ğ4IIk�O!��� ��bx��;��;W ��{�h������MҴ7���ϡ�ϱ�Tm#=��u���A������PV�8`:zc���1���������>��M`x���Ŕ�)=)��'+�*��<+Y�����ռs1�/�SӮs��H��OOZ��\��z�R�&\䚪;|��{W;;d1�3��Q��}9��p8� N��!�׾iy����G�o�u�s���ڀw�������s���=���pi{t�ny�Ό��R��=�#���p�s���4��R����(�8n?��<gkp?�7J`���;�OQ�� ;ӗ��'�=i����Η?/��d�{�O���^�4���GN޴�6��>��(�����r~^���(�p0��z�]�cg~�����s�֞��>d���������{��������R�{qN����@���#<�ӷz��q���w��8_�b�� U+��	�Ґ��r�/��j�H?秮r�� G�=�G���|=�iXw,|� )� g�g�<��ֳ��͏;=x�� ��O�{�@��Aޟ֝��$�T�޹�/�q��i�P%ač��w��>��gT�B���O��
N�Ǹ?��W&u�'�A�x�U�Q��qv��h�@jw �Rr����N� �����6+���ו��A��y���FI�l��ޙ'{}�<:o�H��o��\�؊rj-���������v;2�ӭ(*K���u���;�u	|�"c��:߾cÎ��(�<�^Ń��õIǖ9�\��.	̲��8�x�89�M1?8/��'�sXI������U����$}=sN�h�08� ��ZQ�/E���n��q�ҥ,	R��]_j ��A��i��O�gM�ۉ#��wO�O�����ӁM��$���7q� ���&G��($y?"���^��G"�+��,g9�<� Z��O$ׁ�k�~� �݌���:��݃܊�>�K�>���~>¾(��Ѿ�%�B�L��TrO��_g��ᔮ�,[�~�5�'�ԝ<Fͅ�����C���K�G>.fx����J������A'a d��VU�q��~��G�^I�Ld�?N������;W*�2#�ڜ
�����@�M�`�ݧ��$cq⤡~]��Z^�zt����+��:��� (�W����6���M�A�֗�:�Z w��O���y��W�x������ q�U�O�� w� ;�t<�}~�Zws������G^���^:�� �P�N��(�~� �4ӎ~�)A���@�-��=;SA\� _�F8'$� ����;~\��@����/��i #�<R���M!A�S�j@�;�����q�� t��8��aOʇ��zL���e���=�2��+|�G�� ��LĜ|��'�~���� g��O��t��F!��~���F`UN�s��j6�yO�c���Qc���0��?©"[,<�|�ݷ8T;��v�5�����)~m���H\S��Kg��0rp��NPz�㷵!lH���S ~g� Ҁ|�{��qޣ��X�d�dg��5�}�Gl�,D���~���\ظ�����?�~�ι�u8�GL�8<��w/�1����V<���	��
�Ė�[���I�u)�$q���aY� i�`c���u�����<���?^*M���I�.��3����V���,QG���ϔ	����j���/(����w� �f��w���U��HT�z�`g����*��.
����5n���T�[�8��ni�5����ڹ�;j�;J��y#�������;���YL���Z��4�b�, V��Q��D�`�O��OQ��͚(T@�* ��1�*���b ����$�r��{�w#�
���R�(����ޥ@�2Nc9;���Ub����"�1���!:7^��7+�!b�@l�#��A'>��֡�P�b�(��nN�kZۨ�"R�q鞹�<���K�X�7�#�i-�N�+��k�HE��2��je�}��Б�z�1��_��1�:����&༸̙e<r3�u��� �3�eIc�߷�X���l�z�F�O�#�J
�Э�+BA�(rI秧nje�ʸA����b[c1~������S��c���vK}n$?)ϓ��ެ%�;r� ��Mp~}ɝO� �qR}�o�}��0I�M;�>&u�p�z1�֞��5>g