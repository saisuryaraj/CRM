9��=C)$�pj~�[���ˤ_p����*�z����M?�V�3��a+p�w�:�z��� ĝ��+0�1�Κ9V�� �X��c������U���-���Q��u��F�}�U���Q�)�E���O�>����f���T$��@c��֯$�ȿ>�l�pA��T�V���y������� $q����#�j�΁�`LG#� �^���V1��c�?��N�D� 4�v̇�l�����3]�D�j�`-�]@5���h�qj�>j�O�����?�W��}7���<�99�� *�+]5؃k7w����J�W���y��.��M��0���B��I���f���U2Wh���W����mPc�q�2��!�4&��4� eA#�O���r�Qs���Y��+������f��wN.ḧR8���M��;��z{�*�c����6����b-pD� ���G��?i�=���L�����:�L���ҟ������@�U#�F��SǘB�����?�tl�1�]�+���ri�!�"п�r��"O�8_h{G�M!\���j�h�;����x2�~�?�U�<��󏓀��T*,9��>�M�Z��*r� 0�5��\��>�L��:W�/��9��Q}�a���g�^+�&� o��5FVX9�9��l�;X�>%k���̮8��k��g���^�\1r����#����H[��k2�5�6��zK�_h�֭B��C�϶��;�
�k�9���y�������;.�N�׎ָ={Y��E����S,�'� v�+�������p�xS�Ǹ�c>V��C���"����1�� 
��M6F��>s�V4W�ȉ���1��8��<C�4s�ڵž�,���q�w-��ޏ6�r��X.;���Ymǁ����5����Fk��A����7�0c����=��Ǧ^��-��l��BA��:�U��{J��k���bR�he�s��k[W����(-�gPv�=G��ӝBK#�1�>A��X��G\5��E�y��95|�����Í��*,m�� �M}k�m����� B�s�C_�~���:�8��	矔���}�=׆l!K��-.	���i�6��.�0���5D�������Tz���fӕL����8ۂJ�|Kl`�kˢπ>�~��[{�Z�V��+���}+E�QG��ym&�m�`��Zʻ���	{"���Tg�>�=+���SH#�-�X��-��|c�jZM�9I�$� ��{�R��$�����X�{�"�H:�~^}1V����Ү`��?z���������;�NW��aң�V�2#�&#��ҝ��Ƶ��ֵ��R�NO�m�D��2�+e���$}}zu���Fn��t1��K��z�e�nx��Q|8�����K;~ �:d� :�D�1�p��W���[�w�d_4�a~��+�b*`��#���KR���>n�g�H��k�G;�+�*9��)�C�r"<�� 9�i��Gݤ!�c�ץWy9꣊���Hz�a�P��?s�M\1m��e����C�p�z�������T� �S��l���N����NN��z�����}�X�r';��)��1�ɓ�T����� ��G'�T;a����_Jg?7+Ԝ�#�}ߥ5G=ON‰(;O��J��(�����x �=j@�!�`O<�U�>�#�� �b�8Rr*H�P�	oN{b��ni�����q�J���l�v��c�z�q�]O�6"���OJR��ra���w����D�`��u��q��K۠�t���O���r[6ԏ��kA�;w�� !s��C+,@?�� ��{I�\��[֬K�JB�*�)���ҲW�ocg�C�(�1��	�@#��*E1��+C1���zq��)��Jz�zn>V� n{�/?(�i=~qG� �@	�G������zv�1�??�]����@��R�eX���V�v>�����w�v4�>M�p��8�&�l8����&�}�Ҽ�\`,�9^!=�̯�VN