Z�u#��;��ZPTF:�	�UUeS0��i7Hd�i�@�z米e�SЌ8��Xw��E������ۏ�8�<zt���Ҏ9ܻ��>����9S��^@�)��#�늪���̘�c���9lpx5d�~c�����}��b�q;���|�Z@������Ԅ �ϷJQ��%~��ڞ:�G��hW�����z�pO�1�w�"���� W�z�[�?�&1T|��/����������[����~�3����ޘ �����w�O�h��o�L�S��w ��ߥ:7_Jo�/^riF6���O#� ;��͎i���n��;G�zS��?���v��Ԁp9h���=��q� ��ݱ����Xt����#� y��Lg�!�z�߭5��a�e���@����݆i��8��
z��4���!{g�P!��(�t'�� :k}�x��p!�N1ʁ��}j'$K�R0�q��ژ�}р:�Zf� ��v����1�C'�L�pA<v��A� VS�3��Z,&<��S�Y���Te�ˑ!�cu4�Q�-���y�{⫻����C�=i�H������ʠ��x�}i����9̜�^�b��޿)�<G8<�;�ǭ<cx��}h+ד�$�8��ϭ��� dw�I�� ��Y��9��R�	8<n?����E��m��&�Q@��r������ʁ_.�	��Y7W�)�8 I����y3]�]J�{�� =�Ҹ�5�+���ʠ�0�sS��J�͗"B2H�۸�H��~�G�1���$r�2��q��=ꖄ�N��`;��3q���5��[D��a�F�Z����I6� .:������n���dӮaP�G���մY��=[o�!>h��ˌ����-����9��Oӥ\��N�J��į����O��A �2�W�.��R���cvp>![_�ݾ�p89�:��k�ۤ;��9�P��ZK++�@=?�ּ�}6�I��'S�s��RF�'�`�߼oÚC���מ)rw`c�R�`���!�zt���_��M'q��� �{�N}���;�{Pdu����|�w���.���ЄCȑ2_�Wb�VS�7���V=�1�Ú�^^3H6�q�k+̹.O�ÿZ��|�;c�Dq������m����ֵl��<g�j�#�;֥�ʷh[w�2=-7�ҡ�_�x=��rDn�(�ZZM�M�ۧ�D#��I[�<�1�*���N��%�5b7������ �}u�cM"́ϐ:�Ҿ[�uf�?�^����B�;dC���qZ�Z���OX\}�9o�ڨ͌͝���� ?�c��Eg�pڻbp6eN߼st9�fJ͆�xNjܼ��?LV{n�@c��ִ�J+�N㜚	